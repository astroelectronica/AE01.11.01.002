.title KiCad schematic
.include "models/GBU810.spice.txt"
D1 /LINE VCC DI_GBU810
D2 /NEUTRAL VCC DI_GBU810
D3 0 /LINE DI_GBU810
D4 0 /NEUTRAL DI_GBU810
C1 /VC 0 {CBULK}
R1 VCC /VC {RSER_BULK}
R2 VCC 0 {RLOAD}
V1 /LINE /NEUTRAL SINE({VOFFSET} {VPK} {FREQ})
.end
